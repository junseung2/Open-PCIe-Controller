package pcie_tl_env_pkg;

import uvm_pkg::*;
import pcie_tl_stimulus_pkg::*;

`include "pcie_tl_driver.sv"
`include "pcie_tl_monitor.sv"
`include "pcie_tl_agent.sv"
`include "pcie_tl_scoreboard.sv"
`include "pcie_tl_environment.sv"

endpackage