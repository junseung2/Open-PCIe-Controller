package pcie_tl_stimulus_pkg;

import uvm_pkg::*;

`include "pcie_tl_item.sv"
`include "pcie_tl_sequence.sv"

endpackage