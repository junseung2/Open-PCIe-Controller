package pcie_dll_stimulus_pkg;

import uvm_pkg::*;

`include "pcie_dll_item.sv"
`include "pcie_dll_sequence.sv"

endpackage