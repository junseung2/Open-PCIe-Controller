package pcie_dll_env_pkg;

import uvm_pkg::*;
import pcie_dll_stimulus_pkg::*;

`include "pcie_dll_driver.sv"
`include "pcie_dll_monitor.sv"
`include "pcie_dll_agent.sv"
`include "pcie_dll_scoreboard.sv"
`include "pcie_dll_environment.sv"

endpackage