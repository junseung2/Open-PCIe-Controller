package pcie_tl_test_pkg;

import uvm_pkg::*;
import pcie_tl_stimulus_pkg::*;
import pcie_tl_env_pkg::*;

`include "pcie_tl_base_test.sv"

endpackage