package pcie_dll_test_pkg;

import uvm_pkg::*;
import pcie_dll_stimulus_pkg::*;
import pcie_dll_env_pkg::*;

`include "pcie_dll_base_test.sv"

endpackage